`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Aastha V
// 
// Create Date:    19:07:07 07/15/2019 
// Design Name: 
// Module Name:    dist_RAM_block 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dist_RAM_block(
    output [232:0] out1,
    output [232:0] out2,
    input [232:0] din,
    input [3:0] add1,
    input [3:0] add2,
    input we,
    input clk
    );
	 
// specifications : 
//Single-Port and Dual-Port Distributed RAMs
//  Primitive     RAM Size(Depth x Width)     Type        Address Inputs
//1.RAM16X1S      16 x 1                      Single-port  A3, A2, A1, A0
//2.RAM32X1S      32 x 1 							 Single-port  A4, A3, A2, A1, A0
//3.RAM64X1S 		 64 x 1 							 Single-port  A5, A4, A3, A2, A1, A0
//4.RAM16X1D 		 16 x 1 							 Dual-port    A3, A2, A1, A0

//-------choosen the fourth one---------

wire [232:0] temp_out1, temp_out2;

RAM16X1D ram_0(temp_out2[0], temp_out1[0], add1[0], add1[1], add1[2], add1[3], din[0], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_1(temp_out2[1], temp_out1[1], add1[0], add1[1], add1[2], add1[3], din[1], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_2(temp_out2[2], temp_out1[2], add1[0], add1[1], add1[2], add1[3], din[2], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_3(temp_out2[3], temp_out1[3], add1[0], add1[1], add1[2], add1[3], din[3], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_4(temp_out2[4], temp_out1[4], add1[0], add1[1], add1[2], add1[3], din[4], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_5(temp_out2[5], temp_out1[5], add1[0], add1[1], add1[2], add1[3], din[5], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_6(temp_out2[6], temp_out1[6], add1[0], add1[1], add1[2], add1[3], din[6], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_7(temp_out2[7], temp_out1[7], add1[0], add1[1], add1[2], add1[3], din[7], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_8(temp_out2[8], temp_out1[8], add1[0], add1[1], add1[2], add1[3], din[8], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_9(temp_out2[9], temp_out1[9], add1[0], add1[1], add1[2], add1[3], din[9], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_10(temp_out2[10], temp_out1[10], add1[0], add1[1], add1[2], add1[3], din[10], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_11(temp_out2[11], temp_out1[11], add1[0], add1[1], add1[2], add1[3], din[11], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_12(temp_out2[12], temp_out1[12], add1[0], add1[1], add1[2], add1[3], din[12], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_13(temp_out2[13], temp_out1[13], add1[0], add1[1], add1[2], add1[3], din[13], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_14(temp_out2[14], temp_out1[14], add1[0], add1[1], add1[2], add1[3], din[14], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_15(temp_out2[15], temp_out1[15], add1[0], add1[1], add1[2], add1[3], din[15], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_16(temp_out2[16], temp_out1[16], add1[0], add1[1], add1[2], add1[3], din[16], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_17(temp_out2[17], temp_out1[17], add1[0], add1[1], add1[2], add1[3], din[17], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_18(temp_out2[18], temp_out1[18], add1[0], add1[1], add1[2], add1[3], din[18], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_19(temp_out2[19], temp_out1[19], add1[0], add1[1], add1[2], add1[3], din[19], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_20(temp_out2[20], temp_out1[20], add1[0], add1[1], add1[2], add1[3], din[20], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_21(temp_out2[21], temp_out1[21], add1[0], add1[1], add1[2], add1[3], din[21], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_22(temp_out2[22], temp_out1[22], add1[0], add1[1], add1[2], add1[3], din[22], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_23(temp_out2[23], temp_out1[23], add1[0], add1[1], add1[2], add1[3], din[23], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_24(temp_out2[24], temp_out1[24], add1[0], add1[1], add1[2], add1[3], din[24], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_25(temp_out2[25], temp_out1[25], add1[0], add1[1], add1[2], add1[3], din[25], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_26(temp_out2[26], temp_out1[26], add1[0], add1[1], add1[2], add1[3], din[26], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_27(temp_out2[27], temp_out1[27], add1[0], add1[1], add1[2], add1[3], din[27], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_28(temp_out2[28], temp_out1[28], add1[0], add1[1], add1[2], add1[3], din[28], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_29(temp_out2[29], temp_out1[29], add1[0], add1[1], add1[2], add1[3], din[29], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_30(temp_out2[30], temp_out1[30], add1[0], add1[1], add1[2], add1[3], din[30], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_31(temp_out2[31], temp_out1[31], add1[0], add1[1], add1[2], add1[3], din[31], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_32(temp_out2[32], temp_out1[32], add1[0], add1[1], add1[2], add1[3], din[32], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_33(temp_out2[33], temp_out1[33], add1[0], add1[1], add1[2], add1[3], din[33], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_34(temp_out2[34], temp_out1[34], add1[0], add1[1], add1[2], add1[3], din[34], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_35(temp_out2[35], temp_out1[35], add1[0], add1[1], add1[2], add1[3], din[35], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_36(temp_out2[36], temp_out1[36], add1[0], add1[1], add1[2], add1[3], din[36], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_37(temp_out2[37], temp_out1[37], add1[0], add1[1], add1[2], add1[3], din[37], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_38(temp_out2[38], temp_out1[38], add1[0], add1[1], add1[2], add1[3], din[38], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_39(temp_out2[39], temp_out1[39], add1[0], add1[1], add1[2], add1[3], din[39], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_40(temp_out2[40], temp_out1[40], add1[0], add1[1], add1[2], add1[3], din[40], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_41(temp_out2[41], temp_out1[41], add1[0], add1[1], add1[2], add1[3], din[41], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_42(temp_out2[42], temp_out1[42], add1[0], add1[1], add1[2], add1[3], din[42], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_43(temp_out2[43], temp_out1[43], add1[0], add1[1], add1[2], add1[3], din[43], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_44(temp_out2[44], temp_out1[44], add1[0], add1[1], add1[2], add1[3], din[44], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_45(temp_out2[45], temp_out1[45], add1[0], add1[1], add1[2], add1[3], din[45], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_46(temp_out2[46], temp_out1[46], add1[0], add1[1], add1[2], add1[3], din[46], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_47(temp_out2[47], temp_out1[47], add1[0], add1[1], add1[2], add1[3], din[47], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_48(temp_out2[48], temp_out1[48], add1[0], add1[1], add1[2], add1[3], din[48], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_49(temp_out2[49], temp_out1[49], add1[0], add1[1], add1[2], add1[3], din[49], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_50(temp_out2[50], temp_out1[50], add1[0], add1[1], add1[2], add1[3], din[50], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_51(temp_out2[51], temp_out1[51], add1[0], add1[1], add1[2], add1[3], din[51], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_52(temp_out2[52], temp_out1[52], add1[0], add1[1], add1[2], add1[3], din[52], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_53(temp_out2[53], temp_out1[53], add1[0], add1[1], add1[2], add1[3], din[53], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_54(temp_out2[54], temp_out1[54], add1[0], add1[1], add1[2], add1[3], din[54], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_55(temp_out2[55], temp_out1[55], add1[0], add1[1], add1[2], add1[3], din[55], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_56(temp_out2[56], temp_out1[56], add1[0], add1[1], add1[2], add1[3], din[56], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_57(temp_out2[57], temp_out1[57], add1[0], add1[1], add1[2], add1[3], din[57], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_58(temp_out2[58], temp_out1[58], add1[0], add1[1], add1[2], add1[3], din[58], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_59(temp_out2[59], temp_out1[59], add1[0], add1[1], add1[2], add1[3], din[59], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_60(temp_out2[60], temp_out1[60], add1[0], add1[1], add1[2], add1[3], din[60], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_61(temp_out2[61], temp_out1[61], add1[0], add1[1], add1[2], add1[3], din[61], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_62(temp_out2[62], temp_out1[62], add1[0], add1[1], add1[2], add1[3], din[62], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_63(temp_out2[63], temp_out1[63], add1[0], add1[1], add1[2], add1[3], din[63], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_64(temp_out2[64], temp_out1[64], add1[0], add1[1], add1[2], add1[3], din[64], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_65(temp_out2[65], temp_out1[65], add1[0], add1[1], add1[2], add1[3], din[65], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_66(temp_out2[66], temp_out1[66], add1[0], add1[1], add1[2], add1[3], din[66], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_67(temp_out2[67], temp_out1[67], add1[0], add1[1], add1[2], add1[3], din[67], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_68(temp_out2[68], temp_out1[68], add1[0], add1[1], add1[2], add1[3], din[68], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_69(temp_out2[69], temp_out1[69], add1[0], add1[1], add1[2], add1[3], din[69], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_70(temp_out2[70], temp_out1[70], add1[0], add1[1], add1[2], add1[3], din[70], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_71(temp_out2[71], temp_out1[71], add1[0], add1[1], add1[2], add1[3], din[71], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_72(temp_out2[72], temp_out1[72], add1[0], add1[1], add1[2], add1[3], din[72], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_73(temp_out2[73], temp_out1[73], add1[0], add1[1], add1[2], add1[3], din[73], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_74(temp_out2[74], temp_out1[74], add1[0], add1[1], add1[2], add1[3], din[74], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_75(temp_out2[75], temp_out1[75], add1[0], add1[1], add1[2], add1[3], din[75], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_76(temp_out2[76], temp_out1[76], add1[0], add1[1], add1[2], add1[3], din[76], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_77(temp_out2[77], temp_out1[77], add1[0], add1[1], add1[2], add1[3], din[77], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_78(temp_out2[78], temp_out1[78], add1[0], add1[1], add1[2], add1[3], din[78], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_79(temp_out2[79], temp_out1[79], add1[0], add1[1], add1[2], add1[3], din[79], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_80(temp_out2[80], temp_out1[80], add1[0], add1[1], add1[2], add1[3], din[80], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_81(temp_out2[81], temp_out1[81], add1[0], add1[1], add1[2], add1[3], din[81], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_82(temp_out2[82], temp_out1[82], add1[0], add1[1], add1[2], add1[3], din[82], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_83(temp_out2[83], temp_out1[83], add1[0], add1[1], add1[2], add1[3], din[83], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_84(temp_out2[84], temp_out1[84], add1[0], add1[1], add1[2], add1[3], din[84], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_85(temp_out2[85], temp_out1[85], add1[0], add1[1], add1[2], add1[3], din[85], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_86(temp_out2[86], temp_out1[86], add1[0], add1[1], add1[2], add1[3], din[86], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_87(temp_out2[87], temp_out1[87], add1[0], add1[1], add1[2], add1[3], din[87], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_88(temp_out2[88], temp_out1[88], add1[0], add1[1], add1[2], add1[3], din[88], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_89(temp_out2[89], temp_out1[89], add1[0], add1[1], add1[2], add1[3], din[89], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_90(temp_out2[90], temp_out1[90], add1[0], add1[1], add1[2], add1[3], din[90], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_91(temp_out2[91], temp_out1[91], add1[0], add1[1], add1[2], add1[3], din[91], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_92(temp_out2[92], temp_out1[92], add1[0], add1[1], add1[2], add1[3], din[92], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_93(temp_out2[93], temp_out1[93], add1[0], add1[1], add1[2], add1[3], din[93], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_94(temp_out2[94], temp_out1[94], add1[0], add1[1], add1[2], add1[3], din[94], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_95(temp_out2[95], temp_out1[95], add1[0], add1[1], add1[2], add1[3], din[95], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_96(temp_out2[96], temp_out1[96], add1[0], add1[1], add1[2], add1[3], din[96], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_97(temp_out2[97], temp_out1[97], add1[0], add1[1], add1[2], add1[3], din[97], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_98(temp_out2[98], temp_out1[98], add1[0], add1[1], add1[2], add1[3], din[98], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_99(temp_out2[99], temp_out1[99], add1[0], add1[1], add1[2], add1[3], din[99], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_100(temp_out2[100], temp_out1[100], add1[0], add1[1], add1[2], add1[3], din[100], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_101(temp_out2[101], temp_out1[101], add1[0], add1[1], add1[2], add1[3], din[101], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_102(temp_out2[102], temp_out1[102], add1[0], add1[1], add1[2], add1[3], din[102], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_103(temp_out2[103], temp_out1[103], add1[0], add1[1], add1[2], add1[3], din[103], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_104(temp_out2[104], temp_out1[104], add1[0], add1[1], add1[2], add1[3], din[104], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_105(temp_out2[105], temp_out1[105], add1[0], add1[1], add1[2], add1[3], din[105], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_106(temp_out2[106], temp_out1[106], add1[0], add1[1], add1[2], add1[3], din[106], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_107(temp_out2[107], temp_out1[107], add1[0], add1[1], add1[2], add1[3], din[107], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_108(temp_out2[108], temp_out1[108], add1[0], add1[1], add1[2], add1[3], din[108], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_109(temp_out2[109], temp_out1[109], add1[0], add1[1], add1[2], add1[3], din[109], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_110(temp_out2[110], temp_out1[110], add1[0], add1[1], add1[2], add1[3], din[110], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_111(temp_out2[111], temp_out1[111], add1[0], add1[1], add1[2], add1[3], din[111], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_112(temp_out2[112], temp_out1[112], add1[0], add1[1], add1[2], add1[3], din[112], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_113(temp_out2[113], temp_out1[113], add1[0], add1[1], add1[2], add1[3], din[113], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_114(temp_out2[114], temp_out1[114], add1[0], add1[1], add1[2], add1[3], din[114], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_115(temp_out2[115], temp_out1[115], add1[0], add1[1], add1[2], add1[3], din[115], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_116(temp_out2[116], temp_out1[116], add1[0], add1[1], add1[2], add1[3], din[116], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_117(temp_out2[117], temp_out1[117], add1[0], add1[1], add1[2], add1[3], din[117], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_118(temp_out2[118], temp_out1[118], add1[0], add1[1], add1[2], add1[3], din[118], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_119(temp_out2[119], temp_out1[119], add1[0], add1[1], add1[2], add1[3], din[119], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_120(temp_out2[120], temp_out1[120], add1[0], add1[1], add1[2], add1[3], din[120], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_121(temp_out2[121], temp_out1[121], add1[0], add1[1], add1[2], add1[3], din[121], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_122(temp_out2[122], temp_out1[122], add1[0], add1[1], add1[2], add1[3], din[122], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_123(temp_out2[123], temp_out1[123], add1[0], add1[1], add1[2], add1[3], din[123], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_124(temp_out2[124], temp_out1[124], add1[0], add1[1], add1[2], add1[3], din[124], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_125(temp_out2[125], temp_out1[125], add1[0], add1[1], add1[2], add1[3], din[125], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_126(temp_out2[126], temp_out1[126], add1[0], add1[1], add1[2], add1[3], din[126], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_127(temp_out2[127], temp_out1[127], add1[0], add1[1], add1[2], add1[3], din[127], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_128(temp_out2[128], temp_out1[128], add1[0], add1[1], add1[2], add1[3], din[128], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_129(temp_out2[129], temp_out1[129], add1[0], add1[1], add1[2], add1[3], din[129], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_130(temp_out2[130], temp_out1[130], add1[0], add1[1], add1[2], add1[3], din[130], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_131(temp_out2[131], temp_out1[131], add1[0], add1[1], add1[2], add1[3], din[131], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_132(temp_out2[132], temp_out1[132], add1[0], add1[1], add1[2], add1[3], din[132], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_133(temp_out2[133], temp_out1[133], add1[0], add1[1], add1[2], add1[3], din[133], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_134(temp_out2[134], temp_out1[134], add1[0], add1[1], add1[2], add1[3], din[134], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_135(temp_out2[135], temp_out1[135], add1[0], add1[1], add1[2], add1[3], din[135], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_136(temp_out2[136], temp_out1[136], add1[0], add1[1], add1[2], add1[3], din[136], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_137(temp_out2[137], temp_out1[137], add1[0], add1[1], add1[2], add1[3], din[137], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_138(temp_out2[138], temp_out1[138], add1[0], add1[1], add1[2], add1[3], din[138], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_139(temp_out2[139], temp_out1[139], add1[0], add1[1], add1[2], add1[3], din[139], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_140(temp_out2[140], temp_out1[140], add1[0], add1[1], add1[2], add1[3], din[140], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_141(temp_out2[141], temp_out1[141], add1[0], add1[1], add1[2], add1[3], din[141], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_142(temp_out2[142], temp_out1[142], add1[0], add1[1], add1[2], add1[3], din[142], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_143(temp_out2[143], temp_out1[143], add1[0], add1[1], add1[2], add1[3], din[143], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_144(temp_out2[144], temp_out1[144], add1[0], add1[1], add1[2], add1[3], din[144], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_145(temp_out2[145], temp_out1[145], add1[0], add1[1], add1[2], add1[3], din[145], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_146(temp_out2[146], temp_out1[146], add1[0], add1[1], add1[2], add1[3], din[146], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_147(temp_out2[147], temp_out1[147], add1[0], add1[1], add1[2], add1[3], din[147], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_148(temp_out2[148], temp_out1[148], add1[0], add1[1], add1[2], add1[3], din[148], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_149(temp_out2[149], temp_out1[149], add1[0], add1[1], add1[2], add1[3], din[149], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_150(temp_out2[150], temp_out1[150], add1[0], add1[1], add1[2], add1[3], din[150], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_151(temp_out2[151], temp_out1[151], add1[0], add1[1], add1[2], add1[3], din[151], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_152(temp_out2[152], temp_out1[152], add1[0], add1[1], add1[2], add1[3], din[152], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_153(temp_out2[153], temp_out1[153], add1[0], add1[1], add1[2], add1[3], din[153], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_154(temp_out2[154], temp_out1[154], add1[0], add1[1], add1[2], add1[3], din[154], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_155(temp_out2[155], temp_out1[155], add1[0], add1[1], add1[2], add1[3], din[155], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_156(temp_out2[156], temp_out1[156], add1[0], add1[1], add1[2], add1[3], din[156], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_157(temp_out2[157], temp_out1[157], add1[0], add1[1], add1[2], add1[3], din[157], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_158(temp_out2[158], temp_out1[158], add1[0], add1[1], add1[2], add1[3], din[158], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_159(temp_out2[159], temp_out1[159], add1[0], add1[1], add1[2], add1[3], din[159], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_160(temp_out2[160], temp_out1[160], add1[0], add1[1], add1[2], add1[3], din[160], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_161(temp_out2[161], temp_out1[161], add1[0], add1[1], add1[2], add1[3], din[161], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_162(temp_out2[162], temp_out1[162], add1[0], add1[1], add1[2], add1[3], din[162], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_163(temp_out2[163], temp_out1[163], add1[0], add1[1], add1[2], add1[3], din[163], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_164(temp_out2[164], temp_out1[164], add1[0], add1[1], add1[2], add1[3], din[164], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_165(temp_out2[165], temp_out1[165], add1[0], add1[1], add1[2], add1[3], din[165], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_166(temp_out2[166], temp_out1[166], add1[0], add1[1], add1[2], add1[3], din[166], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_167(temp_out2[167], temp_out1[167], add1[0], add1[1], add1[2], add1[3], din[167], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_168(temp_out2[168], temp_out1[168], add1[0], add1[1], add1[2], add1[3], din[168], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_169(temp_out2[169], temp_out1[169], add1[0], add1[1], add1[2], add1[3], din[169], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_170(temp_out2[170], temp_out1[170], add1[0], add1[1], add1[2], add1[3], din[170], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_171(temp_out2[171], temp_out1[171], add1[0], add1[1], add1[2], add1[3], din[171], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_172(temp_out2[172], temp_out1[172], add1[0], add1[1], add1[2], add1[3], din[172], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_173(temp_out2[173], temp_out1[173], add1[0], add1[1], add1[2], add1[3], din[173], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_174(temp_out2[174], temp_out1[174], add1[0], add1[1], add1[2], add1[3], din[174], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_175(temp_out2[175], temp_out1[175], add1[0], add1[1], add1[2], add1[3], din[175], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_176(temp_out2[176], temp_out1[176], add1[0], add1[1], add1[2], add1[3], din[176], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_177(temp_out2[177], temp_out1[177], add1[0], add1[1], add1[2], add1[3], din[177], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_178(temp_out2[178], temp_out1[178], add1[0], add1[1], add1[2], add1[3], din[178], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_179(temp_out2[179], temp_out1[179], add1[0], add1[1], add1[2], add1[3], din[179], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_180(temp_out2[180], temp_out1[180], add1[0], add1[1], add1[2], add1[3], din[180], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_181(temp_out2[181], temp_out1[181], add1[0], add1[1], add1[2], add1[3], din[181], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_182(temp_out2[182], temp_out1[182], add1[0], add1[1], add1[2], add1[3], din[182], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_183(temp_out2[183], temp_out1[183], add1[0], add1[1], add1[2], add1[3], din[183], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_184(temp_out2[184], temp_out1[184], add1[0], add1[1], add1[2], add1[3], din[184], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_185(temp_out2[185], temp_out1[185], add1[0], add1[1], add1[2], add1[3], din[185], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_186(temp_out2[186], temp_out1[186], add1[0], add1[1], add1[2], add1[3], din[186], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_187(temp_out2[187], temp_out1[187], add1[0], add1[1], add1[2], add1[3], din[187], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_188(temp_out2[188], temp_out1[188], add1[0], add1[1], add1[2], add1[3], din[188], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_189(temp_out2[189], temp_out1[189], add1[0], add1[1], add1[2], add1[3], din[189], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_190(temp_out2[190], temp_out1[190], add1[0], add1[1], add1[2], add1[3], din[190], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_191(temp_out2[191], temp_out1[191], add1[0], add1[1], add1[2], add1[3], din[191], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_192(temp_out2[192], temp_out1[192], add1[0], add1[1], add1[2], add1[3], din[192], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_193(temp_out2[193], temp_out1[193], add1[0], add1[1], add1[2], add1[3], din[193], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_194(temp_out2[194], temp_out1[194], add1[0], add1[1], add1[2], add1[3], din[194], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_195(temp_out2[195], temp_out1[195], add1[0], add1[1], add1[2], add1[3], din[195], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_196(temp_out2[196], temp_out1[196], add1[0], add1[1], add1[2], add1[3], din[196], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_197(temp_out2[197], temp_out1[197], add1[0], add1[1], add1[2], add1[3], din[197], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_198(temp_out2[198], temp_out1[198], add1[0], add1[1], add1[2], add1[3], din[198], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_199(temp_out2[199], temp_out1[199], add1[0], add1[1], add1[2], add1[3], din[199], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_200(temp_out2[200], temp_out1[200], add1[0], add1[1], add1[2], add1[3], din[200], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_201(temp_out2[201], temp_out1[201], add1[0], add1[1], add1[2], add1[3], din[201], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_202(temp_out2[202], temp_out1[202], add1[0], add1[1], add1[2], add1[3], din[202], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_203(temp_out2[203], temp_out1[203], add1[0], add1[1], add1[2], add1[3], din[203], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_204(temp_out2[204], temp_out1[204], add1[0], add1[1], add1[2], add1[3], din[204], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_205(temp_out2[205], temp_out1[205], add1[0], add1[1], add1[2], add1[3], din[205], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_206(temp_out2[206], temp_out1[206], add1[0], add1[1], add1[2], add1[3], din[206], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_207(temp_out2[207], temp_out1[207], add1[0], add1[1], add1[2], add1[3], din[207], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_208(temp_out2[208], temp_out1[208], add1[0], add1[1], add1[2], add1[3], din[208], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_209(temp_out2[209], temp_out1[209], add1[0], add1[1], add1[2], add1[3], din[209], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_210(temp_out2[210], temp_out1[210], add1[0], add1[1], add1[2], add1[3], din[210], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_211(temp_out2[211], temp_out1[211], add1[0], add1[1], add1[2], add1[3], din[211], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_212(temp_out2[212], temp_out1[212], add1[0], add1[1], add1[2], add1[3], din[212], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_213(temp_out2[213], temp_out1[213], add1[0], add1[1], add1[2], add1[3], din[213], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_214(temp_out2[214], temp_out1[214], add1[0], add1[1], add1[2], add1[3], din[214], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_215(temp_out2[215], temp_out1[215], add1[0], add1[1], add1[2], add1[3], din[215], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_216(temp_out2[216], temp_out1[216], add1[0], add1[1], add1[2], add1[3], din[216], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_217(temp_out2[217], temp_out1[217], add1[0], add1[1], add1[2], add1[3], din[217], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_218(temp_out2[218], temp_out1[218], add1[0], add1[1], add1[2], add1[3], din[218], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_219(temp_out2[219], temp_out1[219], add1[0], add1[1], add1[2], add1[3], din[219], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_220(temp_out2[220], temp_out1[220], add1[0], add1[1], add1[2], add1[3], din[220], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_221(temp_out2[221], temp_out1[221], add1[0], add1[1], add1[2], add1[3], din[221], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_222(temp_out2[222], temp_out1[222], add1[0], add1[1], add1[2], add1[3], din[222], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_223(temp_out2[223], temp_out1[223], add1[0], add1[1], add1[2], add1[3], din[223], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_224(temp_out2[224], temp_out1[224], add1[0], add1[1], add1[2], add1[3], din[224], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_225(temp_out2[225], temp_out1[225], add1[0], add1[1], add1[2], add1[3], din[225], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_226(temp_out2[226], temp_out1[226], add1[0], add1[1], add1[2], add1[3], din[226], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_227(temp_out2[227], temp_out1[227], add1[0], add1[1], add1[2], add1[3], din[227], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_228(temp_out2[228], temp_out1[228], add1[0], add1[1], add1[2], add1[3], din[228], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_229(temp_out2[229], temp_out1[229], add1[0], add1[1], add1[2], add1[3], din[229], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_230(temp_out2[230], temp_out1[230], add1[0], add1[1], add1[2], add1[3], din[230], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_231(temp_out2[231], temp_out1[231], add1[0], add1[1], add1[2], add1[3], din[231], add2[0], add2[1], add2[2], add2[3], clk, we);
RAM16X1D ram_232(temp_out2[232], temp_out1[232], add1[0], add1[1], add1[2], add1[3], din[232], add2[0], add2[1], add2[2], add2[3], clk, we);

assign dout1[232:0] = temp_out1[232:0];
assign dout2[232:0] = temp_out2[232:0];

endmodule
